module ADPCM_LUT_ROM(
	input wire [11:0] ADDR,
	output wire [15:0] DATA
);


assign DATA =  (ADDR==12'h000) ? 16'h0002 :
					(ADDR==12'h001) ? 16'h0006 :
					(ADDR==12'h002) ? 16'h000a :
					(ADDR==12'h003) ? 16'h000e :
					(ADDR==12'h004) ? 16'h0012 :
					(ADDR==12'h005) ? 16'h0016 :
					(ADDR==12'h006) ? 16'h001a :
					(ADDR==12'h007) ? 16'h001e :
					(ADDR==12'h008) ? 16'hfffe :
					(ADDR==12'h009) ? 16'hfffa :
					(ADDR==12'h00a) ? 16'hfff6 :
					(ADDR==12'h00b) ? 16'hfff2 :
					(ADDR==12'h00c) ? 16'hffee :
					(ADDR==12'h00d) ? 16'hffea :
					(ADDR==12'h00e) ? 16'hffe6 :
					(ADDR==12'h00f) ? 16'hffe2 :
					(ADDR==12'h010) ? 16'h0002 :
					(ADDR==12'h011) ? 16'h0006 :
					(ADDR==12'h012) ? 16'h000a :
					(ADDR==12'h013) ? 16'h000e :
					(ADDR==12'h014) ? 16'h0013 :
					(ADDR==12'h015) ? 16'h0017 :
					(ADDR==12'h016) ? 16'h001b :
					(ADDR==12'h017) ? 16'h001f :
					(ADDR==12'h018) ? 16'hfffe :
					(ADDR==12'h019) ? 16'hfffa :
					(ADDR==12'h01a) ? 16'hfff6 :
					(ADDR==12'h01b) ? 16'hfff2 :
					(ADDR==12'h01c) ? 16'hffed :
					(ADDR==12'h01d) ? 16'hffe9 :
					(ADDR==12'h01e) ? 16'hffe5 :
					(ADDR==12'h01f) ? 16'hffe1 :
					(ADDR==12'h020) ? 16'h0002 :
					(ADDR==12'h021) ? 16'h0006 :
					(ADDR==12'h022) ? 16'h000b :
					(ADDR==12'h023) ? 16'h000f :
					(ADDR==12'h024) ? 16'h0015 :
					(ADDR==12'h025) ? 16'h0019 :
					(ADDR==12'h026) ? 16'h001e :
					(ADDR==12'h027) ? 16'h0022 :
					(ADDR==12'h028) ? 16'hfffe :
					(ADDR==12'h029) ? 16'hfffa :
					(ADDR==12'h02a) ? 16'hfff5 :
					(ADDR==12'h02b) ? 16'hfff1 :
					(ADDR==12'h02c) ? 16'hffeb :
					(ADDR==12'h02d) ? 16'hffe7 :
					(ADDR==12'h02e) ? 16'hffe2 :
					(ADDR==12'h02f) ? 16'hffde :
					(ADDR==12'h030) ? 16'h0002 :
					(ADDR==12'h031) ? 16'h0007 :
					(ADDR==12'h032) ? 16'h000c :
					(ADDR==12'h033) ? 16'h0011 :
					(ADDR==12'h034) ? 16'h0017 :
					(ADDR==12'h035) ? 16'h001c :
					(ADDR==12'h036) ? 16'h0021 :
					(ADDR==12'h037) ? 16'h0026 :
					(ADDR==12'h038) ? 16'hfffe :
					(ADDR==12'h039) ? 16'hfff9 :
					(ADDR==12'h03a) ? 16'hfff4 :
					(ADDR==12'h03b) ? 16'hffef :
					(ADDR==12'h03c) ? 16'hffe9 :
					(ADDR==12'h03d) ? 16'hffe4 :
					(ADDR==12'h03e) ? 16'hffdf :
					(ADDR==12'h03f) ? 16'hffda :
					(ADDR==12'h040) ? 16'h0002 :
					(ADDR==12'h041) ? 16'h0007 :
					(ADDR==12'h042) ? 16'h000d :
					(ADDR==12'h043) ? 16'h0012 :
					(ADDR==12'h044) ? 16'h0019 :
					(ADDR==12'h045) ? 16'h001e :
					(ADDR==12'h046) ? 16'h0024 :
					(ADDR==12'h047) ? 16'h0029 :
					(ADDR==12'h048) ? 16'hfffe :
					(ADDR==12'h049) ? 16'hfff9 :
					(ADDR==12'h04a) ? 16'hfff3 :
					(ADDR==12'h04b) ? 16'hffee :
					(ADDR==12'h04c) ? 16'hffe7 :
					(ADDR==12'h04d) ? 16'hffe2 :
					(ADDR==12'h04e) ? 16'hffdc :
					(ADDR==12'h04f) ? 16'hffd7 :
					(ADDR==12'h050) ? 16'h0003 :
					(ADDR==12'h051) ? 16'h0009 :
					(ADDR==12'h052) ? 16'h000f :
					(ADDR==12'h053) ? 16'h0015 :
					(ADDR==12'h054) ? 16'h001c :
					(ADDR==12'h055) ? 16'h0022 :
					(ADDR==12'h056) ? 16'h0028 :
					(ADDR==12'h057) ? 16'h002e :
					(ADDR==12'h058) ? 16'hfffd :
					(ADDR==12'h059) ? 16'hfff7 :
					(ADDR==12'h05a) ? 16'hfff1 :
					(ADDR==12'h05b) ? 16'hffeb :
					(ADDR==12'h05c) ? 16'hffe4 :
					(ADDR==12'h05d) ? 16'hffde :
					(ADDR==12'h05e) ? 16'hffd8 :
					(ADDR==12'h05f) ? 16'hffd2 :
					(ADDR==12'h060) ? 16'h0003 :
					(ADDR==12'h061) ? 16'h000a :
					(ADDR==12'h062) ? 16'h0011 :
					(ADDR==12'h063) ? 16'h0018 :
					(ADDR==12'h064) ? 16'h001f :
					(ADDR==12'h065) ? 16'h0026 :
					(ADDR==12'h066) ? 16'h002d :
					(ADDR==12'h067) ? 16'h0034 :
					(ADDR==12'h068) ? 16'hfffd :
					(ADDR==12'h069) ? 16'hfff6 :
					(ADDR==12'h06a) ? 16'hffef :
					(ADDR==12'h06b) ? 16'hffe8 :
					(ADDR==12'h06c) ? 16'hffe1 :
					(ADDR==12'h06d) ? 16'hffda :
					(ADDR==12'h06e) ? 16'hffd3 :
					(ADDR==12'h06f) ? 16'hffcc :
					(ADDR==12'h070) ? 16'h0003 :
					(ADDR==12'h071) ? 16'h000a :
					(ADDR==12'h072) ? 16'h0012 :
					(ADDR==12'h073) ? 16'h0019 :
					(ADDR==12'h074) ? 16'h0022 :
					(ADDR==12'h075) ? 16'h0029 :
					(ADDR==12'h076) ? 16'h0031 :
					(ADDR==12'h077) ? 16'h0038 :
					(ADDR==12'h078) ? 16'hfffd :
					(ADDR==12'h079) ? 16'hfff6 :
					(ADDR==12'h07a) ? 16'hffee :
					(ADDR==12'h07b) ? 16'hffe7 :
					(ADDR==12'h07c) ? 16'hffde :
					(ADDR==12'h07d) ? 16'hffd7 :
					(ADDR==12'h07e) ? 16'hffcf :
					(ADDR==12'h07f) ? 16'hffc8 :
					(ADDR==12'h080) ? 16'h0004 :
					(ADDR==12'h081) ? 16'h000c :
					(ADDR==12'h082) ? 16'h0015 :
					(ADDR==12'h083) ? 16'h001d :
					(ADDR==12'h084) ? 16'h0026 :
					(ADDR==12'h085) ? 16'h002e :
					(ADDR==12'h086) ? 16'h0037 :
					(ADDR==12'h087) ? 16'h003f :
					(ADDR==12'h088) ? 16'hfffc :
					(ADDR==12'h089) ? 16'hfff4 :
					(ADDR==12'h08a) ? 16'hffeb :
					(ADDR==12'h08b) ? 16'hffe3 :
					(ADDR==12'h08c) ? 16'hffda :
					(ADDR==12'h08d) ? 16'hffd2 :
					(ADDR==12'h08e) ? 16'hffc9 :
					(ADDR==12'h08f) ? 16'hffc1 :
					(ADDR==12'h090) ? 16'h0004 :
					(ADDR==12'h091) ? 16'h000d :
					(ADDR==12'h092) ? 16'h0016 :
					(ADDR==12'h093) ? 16'h001f :
					(ADDR==12'h094) ? 16'h0029 :
					(ADDR==12'h095) ? 16'h0032 :
					(ADDR==12'h096) ? 16'h003b :
					(ADDR==12'h097) ? 16'h0044 :
					(ADDR==12'h098) ? 16'hfffc :
					(ADDR==12'h099) ? 16'hfff3 :
					(ADDR==12'h09a) ? 16'hffea :
					(ADDR==12'h09b) ? 16'hffe1 :
					(ADDR==12'h09c) ? 16'hffd7 :
					(ADDR==12'h09d) ? 16'hffce :
					(ADDR==12'h09e) ? 16'hffc5 :
					(ADDR==12'h09f) ? 16'hffbc :
					(ADDR==12'h0a0) ? 16'h0005 :
					(ADDR==12'h0a1) ? 16'h000f :
					(ADDR==12'h0a2) ? 16'h0019 :
					(ADDR==12'h0a3) ? 16'h0023 :
					(ADDR==12'h0a4) ? 16'h002e :
					(ADDR==12'h0a5) ? 16'h0038 :
					(ADDR==12'h0a6) ? 16'h0042 :
					(ADDR==12'h0a7) ? 16'h004c :
					(ADDR==12'h0a8) ? 16'hfffb :
					(ADDR==12'h0a9) ? 16'hfff1 :
					(ADDR==12'h0aa) ? 16'hffe7 :
					(ADDR==12'h0ab) ? 16'hffdd :
					(ADDR==12'h0ac) ? 16'hffd2 :
					(ADDR==12'h0ad) ? 16'hffc8 :
					(ADDR==12'h0ae) ? 16'hffbe :
					(ADDR==12'h0af) ? 16'hffb4 :
					(ADDR==12'h0b0) ? 16'h0005 :
					(ADDR==12'h0b1) ? 16'h0010 :
					(ADDR==12'h0b2) ? 16'h001b :
					(ADDR==12'h0b3) ? 16'h0026 :
					(ADDR==12'h0b4) ? 16'h0032 :
					(ADDR==12'h0b5) ? 16'h003d :
					(ADDR==12'h0b6) ? 16'h0048 :
					(ADDR==12'h0b7) ? 16'h0053 :
					(ADDR==12'h0b8) ? 16'hfffb :
					(ADDR==12'h0b9) ? 16'hfff0 :
					(ADDR==12'h0ba) ? 16'hffe5 :
					(ADDR==12'h0bb) ? 16'hffda :
					(ADDR==12'h0bc) ? 16'hffce :
					(ADDR==12'h0bd) ? 16'hffc3 :
					(ADDR==12'h0be) ? 16'hffb8 :
					(ADDR==12'h0bf) ? 16'hffad :
					(ADDR==12'h0c0) ? 16'h0006 :
					(ADDR==12'h0c1) ? 16'h0012 :
					(ADDR==12'h0c2) ? 16'h001f :
					(ADDR==12'h0c3) ? 16'h002b :
					(ADDR==12'h0c4) ? 16'h0038 :
					(ADDR==12'h0c5) ? 16'h0044 :
					(ADDR==12'h0c6) ? 16'h0051 :
					(ADDR==12'h0c7) ? 16'h005d :
					(ADDR==12'h0c8) ? 16'hfffa :
					(ADDR==12'h0c9) ? 16'hffee :
					(ADDR==12'h0ca) ? 16'hffe1 :
					(ADDR==12'h0cb) ? 16'hffd5 :
					(ADDR==12'h0cc) ? 16'hffc8 :
					(ADDR==12'h0cd) ? 16'hffbc :
					(ADDR==12'h0ce) ? 16'hffaf :
					(ADDR==12'h0cf) ? 16'hffa3 :
					(ADDR==12'h0d0) ? 16'h0006 :
					(ADDR==12'h0d1) ? 16'h0013 :
					(ADDR==12'h0d2) ? 16'h0021 :
					(ADDR==12'h0d3) ? 16'h002e :
					(ADDR==12'h0d4) ? 16'h003d :
					(ADDR==12'h0d5) ? 16'h004a :
					(ADDR==12'h0d6) ? 16'h0058 :
					(ADDR==12'h0d7) ? 16'h0065 :
					(ADDR==12'h0d8) ? 16'hfffa :
					(ADDR==12'h0d9) ? 16'hffed :
					(ADDR==12'h0da) ? 16'hffdf :
					(ADDR==12'h0db) ? 16'hffd2 :
					(ADDR==12'h0dc) ? 16'hffc3 :
					(ADDR==12'h0dd) ? 16'hffb6 :
					(ADDR==12'h0de) ? 16'hffa8 :
					(ADDR==12'h0df) ? 16'hff9b :
					(ADDR==12'h0e0) ? 16'h0007 :
					(ADDR==12'h0e1) ? 16'h0016 :
					(ADDR==12'h0e2) ? 16'h0025 :
					(ADDR==12'h0e3) ? 16'h0034 :
					(ADDR==12'h0e4) ? 16'h0043 :
					(ADDR==12'h0e5) ? 16'h0052 :
					(ADDR==12'h0e6) ? 16'h0061 :
					(ADDR==12'h0e7) ? 16'h0070 :
					(ADDR==12'h0e8) ? 16'hfff9 :
					(ADDR==12'h0e9) ? 16'hffea :
					(ADDR==12'h0ea) ? 16'hffdb :
					(ADDR==12'h0eb) ? 16'hffcc :
					(ADDR==12'h0ec) ? 16'hffbd :
					(ADDR==12'h0ed) ? 16'hffae :
					(ADDR==12'h0ee) ? 16'hff9f :
					(ADDR==12'h0ef) ? 16'hff90 :
					(ADDR==12'h0f0) ? 16'h0008 :
					(ADDR==12'h0f1) ? 16'h0018 :
					(ADDR==12'h0f2) ? 16'h0029 :
					(ADDR==12'h0f3) ? 16'h0039 :
					(ADDR==12'h0f4) ? 16'h004a :
					(ADDR==12'h0f5) ? 16'h005a :
					(ADDR==12'h0f6) ? 16'h006b :
					(ADDR==12'h0f7) ? 16'h007b :
					(ADDR==12'h0f8) ? 16'hfff8 :
					(ADDR==12'h0f9) ? 16'hffe8 :
					(ADDR==12'h0fa) ? 16'hffd7 :
					(ADDR==12'h0fb) ? 16'hffc7 :
					(ADDR==12'h0fc) ? 16'hffb6 :
					(ADDR==12'h0fd) ? 16'hffa6 :
					(ADDR==12'h0fe) ? 16'hff95 :
					(ADDR==12'h0ff) ? 16'hff85 :
					(ADDR==12'h100) ? 16'h0009 :
					(ADDR==12'h101) ? 16'h001b :
					(ADDR==12'h102) ? 16'h002d :
					(ADDR==12'h103) ? 16'h003f :
					(ADDR==12'h104) ? 16'h0052 :
					(ADDR==12'h105) ? 16'h0064 :
					(ADDR==12'h106) ? 16'h0076 :
					(ADDR==12'h107) ? 16'h0088 :
					(ADDR==12'h108) ? 16'hfff7 :
					(ADDR==12'h109) ? 16'hffe5 :
					(ADDR==12'h10a) ? 16'hffd3 :
					(ADDR==12'h10b) ? 16'hffc1 :
					(ADDR==12'h10c) ? 16'hffae :
					(ADDR==12'h10d) ? 16'hff9c :
					(ADDR==12'h10e) ? 16'hff8a :
					(ADDR==12'h10f) ? 16'hff78 :
					(ADDR==12'h110) ? 16'h000a :
					(ADDR==12'h111) ? 16'h001e :
					(ADDR==12'h112) ? 16'h0032 :
					(ADDR==12'h113) ? 16'h0046 :
					(ADDR==12'h114) ? 16'h005a :
					(ADDR==12'h115) ? 16'h006e :
					(ADDR==12'h116) ? 16'h0082 :
					(ADDR==12'h117) ? 16'h0096 :
					(ADDR==12'h118) ? 16'hfff6 :
					(ADDR==12'h119) ? 16'hffe2 :
					(ADDR==12'h11a) ? 16'hffce :
					(ADDR==12'h11b) ? 16'hffba :
					(ADDR==12'h11c) ? 16'hffa6 :
					(ADDR==12'h11d) ? 16'hff92 :
					(ADDR==12'h11e) ? 16'hff7e :
					(ADDR==12'h11f) ? 16'hff6a :
					(ADDR==12'h120) ? 16'h000b :
					(ADDR==12'h121) ? 16'h0021 :
					(ADDR==12'h122) ? 16'h0037 :
					(ADDR==12'h123) ? 16'h004d :
					(ADDR==12'h124) ? 16'h0063 :
					(ADDR==12'h125) ? 16'h0079 :
					(ADDR==12'h126) ? 16'h008f :
					(ADDR==12'h127) ? 16'h00a5 :
					(ADDR==12'h128) ? 16'hfff5 :
					(ADDR==12'h129) ? 16'hffdf :
					(ADDR==12'h12a) ? 16'hffc9 :
					(ADDR==12'h12b) ? 16'hffb3 :
					(ADDR==12'h12c) ? 16'hff9d :
					(ADDR==12'h12d) ? 16'hff87 :
					(ADDR==12'h12e) ? 16'hff71 :
					(ADDR==12'h12f) ? 16'hff5b :
					(ADDR==12'h130) ? 16'h000c :
					(ADDR==12'h131) ? 16'h0024 :
					(ADDR==12'h132) ? 16'h003c :
					(ADDR==12'h133) ? 16'h0054 :
					(ADDR==12'h134) ? 16'h006d :
					(ADDR==12'h135) ? 16'h0085 :
					(ADDR==12'h136) ? 16'h009d :
					(ADDR==12'h137) ? 16'h00b5 :
					(ADDR==12'h138) ? 16'hfff4 :
					(ADDR==12'h139) ? 16'hffdc :
					(ADDR==12'h13a) ? 16'hffc4 :
					(ADDR==12'h13b) ? 16'hffac :
					(ADDR==12'h13c) ? 16'hff93 :
					(ADDR==12'h13d) ? 16'hff7b :
					(ADDR==12'h13e) ? 16'hff63 :
					(ADDR==12'h13f) ? 16'hff4b :
					(ADDR==12'h140) ? 16'h000d :
					(ADDR==12'h141) ? 16'h0027 :
					(ADDR==12'h142) ? 16'h0042 :
					(ADDR==12'h143) ? 16'h005c :
					(ADDR==12'h144) ? 16'h0078 :
					(ADDR==12'h145) ? 16'h0092 :
					(ADDR==12'h146) ? 16'h00ad :
					(ADDR==12'h147) ? 16'h00c7 :
					(ADDR==12'h148) ? 16'hfff3 :
					(ADDR==12'h149) ? 16'hffd9 :
					(ADDR==12'h14a) ? 16'hffbe :
					(ADDR==12'h14b) ? 16'hffa4 :
					(ADDR==12'h14c) ? 16'hff88 :
					(ADDR==12'h14d) ? 16'hff6e :
					(ADDR==12'h14e) ? 16'hff53 :
					(ADDR==12'h14f) ? 16'hff39 :
					(ADDR==12'h150) ? 16'h000e :
					(ADDR==12'h151) ? 16'h002b :
					(ADDR==12'h152) ? 16'h0049 :
					(ADDR==12'h153) ? 16'h0066 :
					(ADDR==12'h154) ? 16'h0084 :
					(ADDR==12'h155) ? 16'h00a1 :
					(ADDR==12'h156) ? 16'h00bf :
					(ADDR==12'h157) ? 16'h00dc :
					(ADDR==12'h158) ? 16'hfff2 :
					(ADDR==12'h159) ? 16'hffd5 :
					(ADDR==12'h15a) ? 16'hffb7 :
					(ADDR==12'h15b) ? 16'hff9a :
					(ADDR==12'h15c) ? 16'hff7c :
					(ADDR==12'h15d) ? 16'hff5f :
					(ADDR==12'h15e) ? 16'hff41 :
					(ADDR==12'h15f) ? 16'hff24 :
					(ADDR==12'h160) ? 16'h0010 :
					(ADDR==12'h161) ? 16'h0030 :
					(ADDR==12'h162) ? 16'h0051 :
					(ADDR==12'h163) ? 16'h0071 :
					(ADDR==12'h164) ? 16'h0092 :
					(ADDR==12'h165) ? 16'h00b2 :
					(ADDR==12'h166) ? 16'h00d3 :
					(ADDR==12'h167) ? 16'h00f3 :
					(ADDR==12'h168) ? 16'hfff0 :
					(ADDR==12'h169) ? 16'hffd0 :
					(ADDR==12'h16a) ? 16'hffaf :
					(ADDR==12'h16b) ? 16'hff8f :
					(ADDR==12'h16c) ? 16'hff6e :
					(ADDR==12'h16d) ? 16'hff4e :
					(ADDR==12'h16e) ? 16'hff2d :
					(ADDR==12'h16f) ? 16'hff0d :
					(ADDR==12'h170) ? 16'h0011 :
					(ADDR==12'h171) ? 16'h0034 :
					(ADDR==12'h172) ? 16'h0058 :
					(ADDR==12'h173) ? 16'h007b :
					(ADDR==12'h174) ? 16'h00a0 :
					(ADDR==12'h175) ? 16'h00c3 :
					(ADDR==12'h176) ? 16'h00e7 :
					(ADDR==12'h177) ? 16'h010a :
					(ADDR==12'h178) ? 16'hffef :
					(ADDR==12'h179) ? 16'hffcc :
					(ADDR==12'h17a) ? 16'hffa8 :
					(ADDR==12'h17b) ? 16'hff85 :
					(ADDR==12'h17c) ? 16'hff60 :
					(ADDR==12'h17d) ? 16'hff3d :
					(ADDR==12'h17e) ? 16'hff19 :
					(ADDR==12'h17f) ? 16'hfef6 :
					(ADDR==12'h180) ? 16'h0013 :
					(ADDR==12'h181) ? 16'h003a :
					(ADDR==12'h182) ? 16'h0061 :
					(ADDR==12'h183) ? 16'h0088 :
					(ADDR==12'h184) ? 16'h00b0 :
					(ADDR==12'h185) ? 16'h00d7 :
					(ADDR==12'h186) ? 16'h00fe :
					(ADDR==12'h187) ? 16'h0125 :
					(ADDR==12'h188) ? 16'hffed :
					(ADDR==12'h189) ? 16'hffc6 :
					(ADDR==12'h18a) ? 16'hff9f :
					(ADDR==12'h18b) ? 16'hff78 :
					(ADDR==12'h18c) ? 16'hff50 :
					(ADDR==12'h18d) ? 16'hff29 :
					(ADDR==12'h18e) ? 16'hff02 :
					(ADDR==12'h18f) ? 16'hfedb :
					(ADDR==12'h190) ? 16'h0015 :
					(ADDR==12'h191) ? 16'h0040 :
					(ADDR==12'h192) ? 16'h006b :
					(ADDR==12'h193) ? 16'h0096 :
					(ADDR==12'h194) ? 16'h00c2 :
					(ADDR==12'h195) ? 16'h00ed :
					(ADDR==12'h196) ? 16'h0118 :
					(ADDR==12'h197) ? 16'h0143 :
					(ADDR==12'h198) ? 16'hffeb :
					(ADDR==12'h199) ? 16'hffc0 :
					(ADDR==12'h19a) ? 16'hff95 :
					(ADDR==12'h19b) ? 16'hff6a :
					(ADDR==12'h19c) ? 16'hff3e :
					(ADDR==12'h19d) ? 16'hff13 :
					(ADDR==12'h19e) ? 16'hfee8 :
					(ADDR==12'h19f) ? 16'hfebd :
					(ADDR==12'h1a0) ? 16'h0017 :
					(ADDR==12'h1a1) ? 16'h0046 :
					(ADDR==12'h1a2) ? 16'h0076 :
					(ADDR==12'h1a3) ? 16'h00a5 :
					(ADDR==12'h1a4) ? 16'h00d5 :
					(ADDR==12'h1a5) ? 16'h0104 :
					(ADDR==12'h1a6) ? 16'h0134 :
					(ADDR==12'h1a7) ? 16'h0163 :
					(ADDR==12'h1a8) ? 16'hffe9 :
					(ADDR==12'h1a9) ? 16'hffba :
					(ADDR==12'h1aa) ? 16'hff8a :
					(ADDR==12'h1ab) ? 16'hff5b :
					(ADDR==12'h1ac) ? 16'hff2b :
					(ADDR==12'h1ad) ? 16'hfefc :
					(ADDR==12'h1ae) ? 16'hfecc :
					(ADDR==12'h1af) ? 16'hfe9d :
					(ADDR==12'h1b0) ? 16'h001a :
					(ADDR==12'h1b1) ? 16'h004e :
					(ADDR==12'h1b2) ? 16'h0082 :
					(ADDR==12'h1b3) ? 16'h00b6 :
					(ADDR==12'h1b4) ? 16'h00eb :
					(ADDR==12'h1b5) ? 16'h011f :
					(ADDR==12'h1b6) ? 16'h0153 :
					(ADDR==12'h1b7) ? 16'h0187 :
					(ADDR==12'h1b8) ? 16'hffe6 :
					(ADDR==12'h1b9) ? 16'hffb2 :
					(ADDR==12'h1ba) ? 16'hff7e :
					(ADDR==12'h1bb) ? 16'hff4a :
					(ADDR==12'h1bc) ? 16'hff15 :
					(ADDR==12'h1bd) ? 16'hfee1 :
					(ADDR==12'h1be) ? 16'hfead :
					(ADDR==12'h1bf) ? 16'hfe79 :
					(ADDR==12'h1c0) ? 16'h001c :
					(ADDR==12'h1c1) ? 16'h0055 :
					(ADDR==12'h1c2) ? 16'h008f :
					(ADDR==12'h1c3) ? 16'h00c8 :
					(ADDR==12'h1c4) ? 16'h0102 :
					(ADDR==12'h1c5) ? 16'h013b :
					(ADDR==12'h1c6) ? 16'h0175 :
					(ADDR==12'h1c7) ? 16'h01ae :
					(ADDR==12'h1c8) ? 16'hffe4 :
					(ADDR==12'h1c9) ? 16'hffab :
					(ADDR==12'h1ca) ? 16'hff71 :
					(ADDR==12'h1cb) ? 16'hff38 :
					(ADDR==12'h1cc) ? 16'hfefe :
					(ADDR==12'h1cd) ? 16'hfec5 :
					(ADDR==12'h1ce) ? 16'hfe8b :
					(ADDR==12'h1cf) ? 16'hfe52 :
					(ADDR==12'h1d0) ? 16'h001f :
					(ADDR==12'h1d1) ? 16'h005e :
					(ADDR==12'h1d2) ? 16'h009d :
					(ADDR==12'h1d3) ? 16'h00dc :
					(ADDR==12'h1d4) ? 16'h011c :
					(ADDR==12'h1d5) ? 16'h015b :
					(ADDR==12'h1d6) ? 16'h019a :
					(ADDR==12'h1d7) ? 16'h01d9 :
					(ADDR==12'h1d8) ? 16'hffe1 :
					(ADDR==12'h1d9) ? 16'hffa2 :
					(ADDR==12'h1da) ? 16'hff63 :
					(ADDR==12'h1db) ? 16'hff24 :
					(ADDR==12'h1dc) ? 16'hfee4 :
					(ADDR==12'h1dd) ? 16'hfea5 :
					(ADDR==12'h1de) ? 16'hfe66 :
					(ADDR==12'h1df) ? 16'hfe27 :
					(ADDR==12'h1e0) ? 16'h0022 :
					(ADDR==12'h1e1) ? 16'h0067 :
					(ADDR==12'h1e2) ? 16'h00ad :
					(ADDR==12'h1e3) ? 16'h00f2 :
					(ADDR==12'h1e4) ? 16'h0139 :
					(ADDR==12'h1e5) ? 16'h017e :
					(ADDR==12'h1e6) ? 16'h01c4 :
					(ADDR==12'h1e7) ? 16'h0209 :
					(ADDR==12'h1e8) ? 16'hffde :
					(ADDR==12'h1e9) ? 16'hff99 :
					(ADDR==12'h1ea) ? 16'hff53 :
					(ADDR==12'h1eb) ? 16'hff0e :
					(ADDR==12'h1ec) ? 16'hfec7 :
					(ADDR==12'h1ed) ? 16'hfe82 :
					(ADDR==12'h1ee) ? 16'hfe3c :
					(ADDR==12'h1ef) ? 16'hfdf7 :
					(ADDR==12'h1f0) ? 16'h0026 :
					(ADDR==12'h1f1) ? 16'h0072 :
					(ADDR==12'h1f2) ? 16'h00bf :
					(ADDR==12'h1f3) ? 16'h010b :
					(ADDR==12'h1f4) ? 16'h0159 :
					(ADDR==12'h1f5) ? 16'h01a5 :
					(ADDR==12'h1f6) ? 16'h01f2 :
					(ADDR==12'h1f7) ? 16'h023e :
					(ADDR==12'h1f8) ? 16'hffda :
					(ADDR==12'h1f9) ? 16'hff8e :
					(ADDR==12'h1fa) ? 16'hff41 :
					(ADDR==12'h1fb) ? 16'hfef5 :
					(ADDR==12'h1fc) ? 16'hfea7 :
					(ADDR==12'h1fd) ? 16'hfe5b :
					(ADDR==12'h1fe) ? 16'hfe0e :
					(ADDR==12'h1ff) ? 16'hfdc2 :
					(ADDR==12'h200) ? 16'h002a :
					(ADDR==12'h201) ? 16'h007e :
					(ADDR==12'h202) ? 16'h00d2 :
					(ADDR==12'h203) ? 16'h0126 :
					(ADDR==12'h204) ? 16'h017b :
					(ADDR==12'h205) ? 16'h01cf :
					(ADDR==12'h206) ? 16'h0223 :
					(ADDR==12'h207) ? 16'h0277 :
					(ADDR==12'h208) ? 16'hffd6 :
					(ADDR==12'h209) ? 16'hff82 :
					(ADDR==12'h20a) ? 16'hff2e :
					(ADDR==12'h20b) ? 16'hfeda :
					(ADDR==12'h20c) ? 16'hfe85 :
					(ADDR==12'h20d) ? 16'hfe31 :
					(ADDR==12'h20e) ? 16'hfddd :
					(ADDR==12'h20f) ? 16'hfd89 :
					(ADDR==12'h210) ? 16'h002e :
					(ADDR==12'h211) ? 16'h008a :
					(ADDR==12'h212) ? 16'h00e7 :
					(ADDR==12'h213) ? 16'h0143 :
					(ADDR==12'h214) ? 16'h01a1 :
					(ADDR==12'h215) ? 16'h01fd :
					(ADDR==12'h216) ? 16'h025a :
					(ADDR==12'h217) ? 16'h02b6 :
					(ADDR==12'h218) ? 16'hffd2 :
					(ADDR==12'h219) ? 16'hff76 :
					(ADDR==12'h21a) ? 16'hff19 :
					(ADDR==12'h21b) ? 16'hfebd :
					(ADDR==12'h21c) ? 16'hfe5f :
					(ADDR==12'h21d) ? 16'hfe03 :
					(ADDR==12'h21e) ? 16'hfda6 :
					(ADDR==12'h21f) ? 16'hfd4a :
					(ADDR==12'h220) ? 16'h0033 :
					(ADDR==12'h221) ? 16'h0099 :
					(ADDR==12'h222) ? 16'h00ff :
					(ADDR==12'h223) ? 16'h0165 :
					(ADDR==12'h224) ? 16'h01cb :
					(ADDR==12'h225) ? 16'h0231 :
					(ADDR==12'h226) ? 16'h0297 :
					(ADDR==12'h227) ? 16'h02fd :
					(ADDR==12'h228) ? 16'hffcd :
					(ADDR==12'h229) ? 16'hff67 :
					(ADDR==12'h22a) ? 16'hff01 :
					(ADDR==12'h22b) ? 16'hfe9b :
					(ADDR==12'h22c) ? 16'hfe35 :
					(ADDR==12'h22d) ? 16'hfdcf :
					(ADDR==12'h22e) ? 16'hfd69 :
					(ADDR==12'h22f) ? 16'hfd03 :
					(ADDR==12'h230) ? 16'h0038 :
					(ADDR==12'h231) ? 16'h00a8 :
					(ADDR==12'h232) ? 16'h0118 :
					(ADDR==12'h233) ? 16'h0188 :
					(ADDR==12'h234) ? 16'h01f9 :
					(ADDR==12'h235) ? 16'h0269 :
					(ADDR==12'h236) ? 16'h02d9 :
					(ADDR==12'h237) ? 16'h0349 :
					(ADDR==12'h238) ? 16'hffc8 :
					(ADDR==12'h239) ? 16'hff58 :
					(ADDR==12'h23a) ? 16'hfee8 :
					(ADDR==12'h23b) ? 16'hfe78 :
					(ADDR==12'h23c) ? 16'hfe07 :
					(ADDR==12'h23d) ? 16'hfd97 :
					(ADDR==12'h23e) ? 16'hfd27 :
					(ADDR==12'h23f) ? 16'hfcb7 :
					(ADDR==12'h240) ? 16'h003d :
					(ADDR==12'h241) ? 16'h00b8 :
					(ADDR==12'h242) ? 16'h0134 :
					(ADDR==12'h243) ? 16'h01af :
					(ADDR==12'h244) ? 16'h022b :
					(ADDR==12'h245) ? 16'h02a6 :
					(ADDR==12'h246) ? 16'h0322 :
					(ADDR==12'h247) ? 16'h039d :
					(ADDR==12'h248) ? 16'hffc3 :
					(ADDR==12'h249) ? 16'hff48 :
					(ADDR==12'h24a) ? 16'hfecc :
					(ADDR==12'h24b) ? 16'hfe51 :
					(ADDR==12'h24c) ? 16'hfdd5 :
					(ADDR==12'h24d) ? 16'hfd5a :
					(ADDR==12'h24e) ? 16'hfcde :
					(ADDR==12'h24f) ? 16'hfc63 :
					(ADDR==12'h250) ? 16'h0044 :
					(ADDR==12'h251) ? 16'h00cc :
					(ADDR==12'h252) ? 16'h0154 :
					(ADDR==12'h253) ? 16'h01dc :
					(ADDR==12'h254) ? 16'h0264 :
					(ADDR==12'h255) ? 16'h02ec :
					(ADDR==12'h256) ? 16'h0374 :
					(ADDR==12'h257) ? 16'h03fc :
					(ADDR==12'h258) ? 16'hffbc :
					(ADDR==12'h259) ? 16'hff34 :
					(ADDR==12'h25a) ? 16'hfeac :
					(ADDR==12'h25b) ? 16'hfe24 :
					(ADDR==12'h25c) ? 16'hfd9c :
					(ADDR==12'h25d) ? 16'hfd14 :
					(ADDR==12'h25e) ? 16'hfc8c :
					(ADDR==12'h25f) ? 16'hfc04 :
					(ADDR==12'h260) ? 16'h004a :
					(ADDR==12'h261) ? 16'h00df :
					(ADDR==12'h262) ? 16'h0175 :
					(ADDR==12'h263) ? 16'h020a :
					(ADDR==12'h264) ? 16'h02a0 :
					(ADDR==12'h265) ? 16'h0335 :
					(ADDR==12'h266) ? 16'h03cb :
					(ADDR==12'h267) ? 16'h0460 :
					(ADDR==12'h268) ? 16'hffb6 :
					(ADDR==12'h269) ? 16'hff21 :
					(ADDR==12'h26a) ? 16'hfe8b :
					(ADDR==12'h26b) ? 16'hfdf6 :
					(ADDR==12'h26c) ? 16'hfd60 :
					(ADDR==12'h26d) ? 16'hfccb :
					(ADDR==12'h26e) ? 16'hfc35 :
					(ADDR==12'h26f) ? 16'hfba0 :
					(ADDR==12'h270) ? 16'h0052 :
					(ADDR==12'h271) ? 16'h00f6 :
					(ADDR==12'h272) ? 16'h019b :
					(ADDR==12'h273) ? 16'h023f :
					(ADDR==12'h274) ? 16'h02e4 :
					(ADDR==12'h275) ? 16'h0388 :
					(ADDR==12'h276) ? 16'h042d :
					(ADDR==12'h277) ? 16'h04d1 :
					(ADDR==12'h278) ? 16'hffae :
					(ADDR==12'h279) ? 16'hff0a :
					(ADDR==12'h27a) ? 16'hfe65 :
					(ADDR==12'h27b) ? 16'hfdc1 :
					(ADDR==12'h27c) ? 16'hfd1c :
					(ADDR==12'h27d) ? 16'hfc78 :
					(ADDR==12'h27e) ? 16'hfbd3 :
					(ADDR==12'h27f) ? 16'hfb2f :
					(ADDR==12'h280) ? 16'h005a :
					(ADDR==12'h281) ? 16'h010f :
					(ADDR==12'h282) ? 16'h01c4 :
					(ADDR==12'h283) ? 16'h0279 :
					(ADDR==12'h284) ? 16'h032e :
					(ADDR==12'h285) ? 16'h03e3 :
					(ADDR==12'h286) ? 16'h0498 :
					(ADDR==12'h287) ? 16'h054d :
					(ADDR==12'h288) ? 16'hffa6 :
					(ADDR==12'h289) ? 16'hfef1 :
					(ADDR==12'h28a) ? 16'hfe3c :
					(ADDR==12'h28b) ? 16'hfd87 :
					(ADDR==12'h28c) ? 16'hfcd2 :
					(ADDR==12'h28d) ? 16'hfc1d :
					(ADDR==12'h28e) ? 16'hfb68 :
					(ADDR==12'h28f) ? 16'hfab3 :
					(ADDR==12'h290) ? 16'h0063 :
					(ADDR==12'h291) ? 16'h012a :
					(ADDR==12'h292) ? 16'h01f1 :
					(ADDR==12'h293) ? 16'h02b8 :
					(ADDR==12'h294) ? 16'h037f :
					(ADDR==12'h295) ? 16'h0446 :
					(ADDR==12'h296) ? 16'h050d :
					(ADDR==12'h297) ? 16'h05d4 :
					(ADDR==12'h298) ? 16'hff9d :
					(ADDR==12'h299) ? 16'hfed6 :
					(ADDR==12'h29a) ? 16'hfe0f :
					(ADDR==12'h29b) ? 16'hfd48 :
					(ADDR==12'h29c) ? 16'hfc81 :
					(ADDR==12'h29d) ? 16'hfbba :
					(ADDR==12'h29e) ? 16'hfaf3 :
					(ADDR==12'h29f) ? 16'hfa2c :
					(ADDR==12'h2a0) ? 16'h006d :
					(ADDR==12'h2a1) ? 16'h0148 :
					(ADDR==12'h2a2) ? 16'h0223 :
					(ADDR==12'h2a3) ? 16'h02fe :
					(ADDR==12'h2a4) ? 16'h03d9 :
					(ADDR==12'h2a5) ? 16'h04b4 :
					(ADDR==12'h2a6) ? 16'h058f :
					(ADDR==12'h2a7) ? 16'h066a :
					(ADDR==12'h2a8) ? 16'hff93 :
					(ADDR==12'h2a9) ? 16'hfeb8 :
					(ADDR==12'h2aa) ? 16'hfddd :
					(ADDR==12'h2ab) ? 16'hfd02 :
					(ADDR==12'h2ac) ? 16'hfc27 :
					(ADDR==12'h2ad) ? 16'hfb4c :
					(ADDR==12'h2ae) ? 16'hfa71 :
					(ADDR==12'h2af) ? 16'hf996 :
					(ADDR==12'h2b0) ? 16'h0078 :
					(ADDR==12'h2b1) ? 16'h0168 :
					(ADDR==12'h2b2) ? 16'h0259 :
					(ADDR==12'h2b3) ? 16'h0349 :
					(ADDR==12'h2b4) ? 16'h043b :
					(ADDR==12'h2b5) ? 16'h052b :
					(ADDR==12'h2b6) ? 16'h061c :
					(ADDR==12'h2b7) ? 16'h070c :
					(ADDR==12'h2b8) ? 16'hff88 :
					(ADDR==12'h2b9) ? 16'hfe98 :
					(ADDR==12'h2ba) ? 16'hfda7 :
					(ADDR==12'h2bb) ? 16'hfcb7 :
					(ADDR==12'h2bc) ? 16'hfbc5 :
					(ADDR==12'h2bd) ? 16'hfad5 :
					(ADDR==12'h2be) ? 16'hf9e4 :
					(ADDR==12'h2bf) ? 16'hf8f4 :
					(ADDR==12'h2c0) ? 16'h0084 :
					(ADDR==12'h2c1) ? 16'h018d :
					(ADDR==12'h2c2) ? 16'h0296 :
					(ADDR==12'h2c3) ? 16'h039f :
					(ADDR==12'h2c4) ? 16'h04a8 :
					(ADDR==12'h2c5) ? 16'h05b1 :
					(ADDR==12'h2c6) ? 16'h06ba :
					(ADDR==12'h2c7) ? 16'h07c3 :
					(ADDR==12'h2c8) ? 16'hff7c :
					(ADDR==12'h2c9) ? 16'hfe73 :
					(ADDR==12'h2ca) ? 16'hfd6a :
					(ADDR==12'h2cb) ? 16'hfc61 :
					(ADDR==12'h2cc) ? 16'hfb58 :
					(ADDR==12'h2cd) ? 16'hfa4f :
					(ADDR==12'h2ce) ? 16'hf946 :
					(ADDR==12'h2cf) ? 16'hf83d :
					(ADDR==12'h2d0) ? 16'h0091 :
					(ADDR==12'h2d1) ? 16'h01b4 :
					(ADDR==12'h2d2) ? 16'h02d8 :
					(ADDR==12'h2d3) ? 16'h03fb :
					(ADDR==12'h2d4) ? 16'h051f :
					(ADDR==12'h2d5) ? 16'h0642 :
					(ADDR==12'h2d6) ? 16'h0766 :
					(ADDR==12'h2d7) ? 16'h0889 :
					(ADDR==12'h2d8) ? 16'hff6f :
					(ADDR==12'h2d9) ? 16'hfe4c :
					(ADDR==12'h2da) ? 16'hfd28 :
					(ADDR==12'h2db) ? 16'hfc05 :
					(ADDR==12'h2dc) ? 16'hfae1 :
					(ADDR==12'h2dd) ? 16'hf9be :
					(ADDR==12'h2de) ? 16'hf89a :
					(ADDR==12'h2df) ? 16'hf777 :
					(ADDR==12'h2e0) ? 16'h00a0 :
					(ADDR==12'h2e1) ? 16'h01e0 :
					(ADDR==12'h2e2) ? 16'h0321 :
					(ADDR==12'h2e3) ? 16'h0461 :
					(ADDR==12'h2e4) ? 16'h05a2 :
					(ADDR==12'h2e5) ? 16'h06e2 :
					(ADDR==12'h2e6) ? 16'h0823 :
					(ADDR==12'h2e7) ? 16'h0963 :
					(ADDR==12'h2e8) ? 16'hff60 :
					(ADDR==12'h2e9) ? 16'hfe20 :
					(ADDR==12'h2ea) ? 16'hfcdf :
					(ADDR==12'h2eb) ? 16'hfb9f :
					(ADDR==12'h2ec) ? 16'hfa5e :
					(ADDR==12'h2ed) ? 16'hf91e :
					(ADDR==12'h2ee) ? 16'hf7dd :
					(ADDR==12'h2ef) ? 16'hf69d :
					(ADDR==12'h2f0) ? 16'h00b0 :
					(ADDR==12'h2f1) ? 16'h0210 :
					(ADDR==12'h2f2) ? 16'h0371 :
					(ADDR==12'h2f3) ? 16'h04d1 :
					(ADDR==12'h2f4) ? 16'h0633 :
					(ADDR==12'h2f5) ? 16'h0793 :
					(ADDR==12'h2f6) ? 16'h08f4 :
					(ADDR==12'h2f7) ? 16'h0a54 :
					(ADDR==12'h2f8) ? 16'hff50 :
					(ADDR==12'h2f9) ? 16'hfdf0 :
					(ADDR==12'h2fa) ? 16'hfc8f :
					(ADDR==12'h2fb) ? 16'hfb2f :
					(ADDR==12'h2fc) ? 16'hf9cd :
					(ADDR==12'h2fd) ? 16'hf86d :
					(ADDR==12'h2fe) ? 16'hf70c :
					(ADDR==12'h2ff) ? 16'hf5ac :
					(ADDR==12'h300) ? 16'h00c2 :
					(ADDR==12'h301) ? 16'h0246 :
					(ADDR==12'h302) ? 16'h03ca :
					(ADDR==12'h303) ? 16'h054e :
					(ADDR==12'h304) ? 16'h06d2 :
					(ADDR==12'h305) ? 16'h0856 :
					(ADDR==12'h306) ? 16'h09da :
					(ADDR==12'h307) ? 16'h0b5e :
					(ADDR==12'h308) ? 16'hff3e :
					(ADDR==12'h309) ? 16'hfdba :
					(ADDR==12'h30a) ? 16'hfc36 :
					(ADDR==12'h30b) ? 16'hfab2 :
					(ADDR==12'h30c) ? 16'hf92e :
					(ADDR==12'h30d) ? 16'hf7aa :
					(ADDR==12'h30e) ? 16'hf626 :
											16'hf4a2;


endmodule
